* Digital Inverter Spice Netlist for ngspice

* Sources
Vin I 0 dc pulse(0 5 100p 1p 1p 100p 200p)
Vdd VDD 0 dc 5

* Main circuit
X1 I ZN VDD VDD 0 0 gf180mcu_fd_sc_mcu7t5v0__inv_1

* Temperature set
.temp 25
.options tnom=25

* Analyses
.control
tran 1p 200p
meas tran high_in FIND V(ZN) AT=100p
meas tran low_in  FIND V(ZN) AT=200p

wrdata inv_simulated.csv {high_in} {low_in}

.endc

* Libraries calling
.include "design.ngspice"
.lib "sm141064.ngspice" typical

.SUBCKT gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
xM_i_0 ZN I VSS VPW nmos_6p0 W=8.2e-07 L=6e-07
xM_i_1 ZN I VDD VNW pmos_6p0 W=1.22e-06 L=5e-07
.ENDS


.end